library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.my.all;

ENTITY SYNC IS
	PORT (
		CLK: IN STD_LOGIC;
		HSYNC, VSYNC: OUT STD_LOGIC;
		R, G, B: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		DATA: IN STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END SYNC;

ARCHITECTURE MAIN OF SYNC IS
	
	SIGNAL RGB: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL HPOS: INTEGER RANGE 0 TO 1688 := 0;
	SIGNAL VPOS: INTEGER RANGE 0 TO 1066 := 0;
	SIGNAL PIXEL: STD_LOGIC;
	SIGNAL PIXEL_ROW: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL PIXEL_COLUMN: STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL ROM_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL NUMBER, POSITION: INTEGER RANGE 0 TO 40 := 0;
	SIGNAL ADDR: STD_LOGIC_VECTOR(6 DOWNTO 0);	
	
	COMPONENT fontROM IS
		PORT(
			clkA: IN STD_LOGIC;
			addrA: IN STD_LOGIC_VECTOR(10 DOWNTO 0);
			dataOutA: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT fontROM;
	
BEGIN
	PROCESS(CLK)
		VARIABLE ANT : INTEGER := 360;	
	BEGIN		
		IF (CLK'EVENT AND CLK = '1') THEN
			IF (HPOS - ANT = 32) THEN
				POSITION <= (POSITION + 1) MOD 40;
				ANT := HPOS;
			END IF;
			IF (HPOS >= 590 AND HPOS <= 720 AND VPOS >= 400 AND VPOS <= 500) THEN
				R <= (OTHERS => PIXEL);
				G <= (OTHERS => PIXEL);
				B <= (OTHERS => PIXEL);
			END IF;

			IF (HPOS < 1688) THEN
				HPOS <= HPOS + 1;
			ELSE
				HPOS <= 0;
				ANT := 360;
				IF (VPOS < 1066) THEN
					VPOS <= VPOS + 1;
				ELSE
					VPOS <= 0;
				END IF;
			END IF;
			
			IF (HPOS > 0	 AND HPOS < 112) THEN
				HSYNC <= '0';
			ELSE
				HSYNC <= '1';
			END IF;
			
			IF (VPOS > 0 AND VPOS < 4) THEN
				VSYNC <= '0';
			ELSE
				VSYNC <= '1';
			END IF;
			
			IF (HPOS >= 0  AND HPOS < 590) OR (VPOS >= 0 AND VPOS <= 400) THEN
				R <= (OTHERS => '0');
				G <= (OTHERS => '0');
				B <= (OTHERS => '0');
			END IF;
			
			IF ((HPOS > 720) OR (VPOS > 500)) THEN
				R <= (OTHERS => '0');
				G <= (OTHERS => '0');
				B <= (OTHERS => '0');
			END IF;
		END IF;
	END PROCESS;
	
	ADDR <= DATA;
	FONT_COMPONENT: fontROM PORT MAP(CLK, ADDR & PIXEL_ROW, ROM_DATA);
	
	PIXEL_ROW <= STD_LOGIC_VECTOR(TO_UNSIGNED(VPOS, 4));
	-- PIXEL_ROW <= STD_LOGIC_VECTOR(TO_UNSIGNED(VPOS, 4))(7 DOWNTO 4);
	PIXEL_COLUMN <= STD_LOGIC_VECTOR(TO_UNSIGNED(HPOS, 3));
	-- PIXEL_COLUMN <= STD_LOGIC_VECTOR(TO_UNSIGNED(HPOS, 3));(7 DOWNTO 4);
	
	PIXEL <= ROM_DATA(7) WHEN PIXEL_COLUMN(2 DOWNTO 0) = "000" ELSE
			ROM_DATA(6) WHEN PIXEL_COLUMN(2 DOWNTO 0) = "001" ELSE
			ROM_DATA(5) WHEN PIXEL_COLUMN(2 DOWNTO 0) = "010" ELSE
			ROM_DATA(4) WHEN PIXEL_COLUMN(2 DOWNTO 0) = "011" ELSE
			ROM_DATA(3) WHEN PIXEL_COLUMN(2 DOWNTO 0) = "100" ELSE
			ROM_DATA(2) WHEN PIXEL_COLUMN(2 DOWNTO 0) = "101" ELSE
			ROM_DATA(1) WHEN PIXEL_COLUMN(2 DOWNTO 0) = "110" ELSE
			ROM_DATA(0) WHEN PIXEL_COLUMN(2 DOWNTO 0) = "111" ELSE '0'; 
	
END MAIN;
		
		
